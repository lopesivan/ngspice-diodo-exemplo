* exemplo de diodo

.include spice_models/D1N4148.mod

vin 1 0 5
r1  1 2 2.5k
d1  2 0 D1N4148

.op
.control
run
print all
.endc
.end
